module full_adder (
input a, 
input b, 
input cin,
output s, 
output cout
);

assign sum = a ^ b ^ cin;
assign cout = (a & b) | (a & cin) | (b & cin);

endmodule